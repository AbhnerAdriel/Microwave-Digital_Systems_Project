module microwave;

endmodule